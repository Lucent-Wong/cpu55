library verilog;
use verilog.vl_types.all;
entity iram_tb is
end iram_tb;
