library verilog;
use verilog.vl_types.all;
entity mux32x32_tb is
end mux32x32_tb;
