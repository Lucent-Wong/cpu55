library verilog;
use verilog.vl_types.all;
entity wfb_tb is
end wfb_tb;
