library verilog;
use verilog.vl_types.all;
entity myreg_tb is
end myreg_tb;
