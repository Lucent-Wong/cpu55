library verilog;
use verilog.vl_types.all;
entity cu_tb is
end cu_tb;
